set object 1 rect from  20 , 100 to 7 , 100 fc rgb "cyan" fillstyle solid
set object 2 rect from 8 , 20 to 7 , 100 fc rgb "cyan" fillstyle solid
set object 3 rect from 4 , 8 to 7 , 100 fc rgb "cyan" fillstyle solid
set object 4 rect from 2 , 4 to 7 , 100 fc rgb "cyan" fillstyle solid
set object 5 rect from 1 , 2 to 7 , 100 fc rgb "cyan" fillstyle solid
set object 6 rect from 0.5 , 1 to 7 , 100 fc rgb "cyan" fillstyle solid
set object 7 rect from 0.25 , 0.5 to 7 , 100 fc rgb "cyan" fillstyle solid
set object 8 rect from 0.18 , 0.25 to 7 , 100 fc rgb "cyan" fillstyle solid
set object 9 rect from 0.15 , 0.18 to 7 , 100 fc rgb "cyan" fillstyle solid
set object 10 rect from 20 , 100 to 5 , 7 fc rgb "cyan" fillstyle solid
set object 11 rect from 8 , 20 to 5 , 7 fc rgb "cyan" fillstyle solid
set object 12 rect from 4 , 8 to 5 , 7 fc rgb "cyan" fillstyle solid
set object 13 rect from 2 , 4 to 5 , 7 fc rgb "cyan" fillstyle solid
set object 14 rect from 1 , 2 to 5 , 7 fc rgb "cyan" fillstyle solid
set object 15 rect from 0.5 , 1 to 5 , 7 fc rgb "cyan" fillstyle solid
set object 16 rect from 0.25 , 0.5 to 5 , 7 fc rgb "cyan" fillstyle solid
set object 17 rect from 0.18 , 0.25 to 5 , 7 fc rgb "cyan" fillstyle solid
set object 18 rect from 0.15 , 0.18 to 5 , 7 fc rgb "cyan" fillstyle solid
set object 19 rect from 20 , 100 to 3 , 5 fc rgb "cyan" fillstyle solid
set object 20 rect from 8 , 20 to 3 , 5 fc rgb "cyan" fillstyle solid
set object 21 rect from 4 , 8 to 3 , 5 fc rgb "cyan" fillstyle solid
set object 22 rect from 2 , 4 to 3 , 5 fc rgb "cyan" fillstyle solid
set object 23 rect from 1 , 2 to 3 , 5 fc rgb "cyan" fillstyle solid
set object 24 rect from 0.5 , 1 to 3 , 5 fc rgb "cyan" fillstyle solid
set object 25 rect from 0.25 , 0.5 to 3 , 5 fc rgb "cyan" fillstyle solid
set object 26 rect from 0.18 , 0.25 to 3 , 5 fc rgb "cyan" fillstyle solid
set object 27 rect from 0.15 , 0.18 to 3 , 5 fc rgb "cyan" fillstyle solid
set object 28 rect from 20 , 100 to 2 , 3 fc rgb "cyan" fillstyle solid
set object 29 rect from 8 , 20 to 2 , 3 fc rgb "cyan" fillstyle solid
set object 30 rect from 4 , 8 to 2 , 3 fc rgb "cyan" fillstyle solid
set object 31 rect from 2 , 4 to 2 , 3 fc rgb "cyan" fillstyle solid
set object 32 rect from 1 , 2 to 2 , 3 fc rgb "cyan" fillstyle solid
set object 33 rect from 0.5 , 1 to 2 , 3 fc rgb "cyan" fillstyle solid
set object 34 rect from 0.25 , 0.5 to 2 , 3 fc rgb "cyan" fillstyle solid
set object 35 rect from 0.18 , 0.25 to 2 , 3 fc rgb "cyan" fillstyle solid
set object 36 rect from 0.15 , 0.18 to 2 , 3 fc rgb "cyan" fillstyle solid
set object 37 rect from 20 , 100 to 1.68 , 2 fc rgb "cyan" fillstyle solid
set object 38 rect from 8 , 20 to 1.68 , 2 fc rgb "cyan" fillstyle solid
set object 39 rect from 4 , 8 to 1.68 , 2 fc rgb "cyan" fillstyle solid
set object 40 rect from 2 , 4 to 1.68 , 2 fc rgb "cyan" fillstyle solid
set object 41 rect from 1 , 2 to 1.68 , 2 fc rgb "cyan" fillstyle solid
set object 42 rect from 0.5 , 1 to 1.68 , 2 fc rgb "cyan" fillstyle solid
set object 43 rect from 0.25 , 0.5 to 1.68 , 2 fc rgb "cyan" fillstyle solid
set object 44 rect from 0.18 , 0.25 to 1.68 , 2 fc rgb "cyan" fillstyle solid
set object 45 rect from 0.15 , 0.18 to 1.68 , 2 fc rgb "cyan" fillstyle solid
set object 46 rect from 20 , 100 to 1.26 , 1.68 fc rgb "cyan" fillstyle solid
set object 47 rect from 8 , 20 to 1.26 , 1.68 fc rgb "cyan" fillstyle solid
set object 48 rect from 4 , 8 to 1.26 , 1.68 fc rgb "cyan" fillstyle solid
set object 49 rect from 2 , 4 to 1.26 , 1.68 fc rgb "cyan" fillstyle solid
set object 50 rect from 1 , 2 to 1.26 , 1.68 fc rgb "cyan" fillstyle solid
set object 51 rect from 0.5 , 1 to 1.26 , 1.68 fc rgb "cyan" fillstyle solid
set object 52 rect from 0.25 , 0.5 to 1.26 , 1.68 fc rgb "cyan" fillstyle solid
set object 53 rect from 0.18 , 0.25 to 1.26 , 1.68 fc rgb "cyan" fillstyle solid
set object 54 rect from 0.15 , 0.18 to 1.26 , 1.68 fc rgb "cyan" fillstyle solid
set object 55 rect from 20 , 100 to 1 , 1.26 fc rgb "cyan" fillstyle solid
set object 56 rect from 8 , 20 to 1 , 1.26 fc rgb "cyan" fillstyle solid
set object 57 rect from 4 , 8 to 1 , 1.26 fc rgb "cyan" fillstyle solid
set object 58 rect from 2 , 4 to 1 , 1.26 fc rgb "cyan" fillstyle solid
set object 59 rect from 1 , 2 to 1 , 1.26 fc rgb "cyan" fillstyle solid
set object 60 rect from 0.5 , 1 to 1 , 1.26 fc rgb "cyan" fillstyle solid
set object 61 rect from 0.25 , 0.5 to 1 , 1.26 fc rgb "cyan" fillstyle solid
set object 62 rect from 0.18 , 0.25 to 1 , 1.26 fc rgb "cyan" fillstyle solid
set object 63 rect from 0.15 , 0.18 to 1 , 1.26 fc rgb "cyan" fillstyle solid
set object 64 rect from 20 , 100 to 0.84 , 1 fc rgb "cyan" fillstyle solid
set object 65 rect from 8 , 20 to 0.84 , 1 fc rgb "cyan" fillstyle solid
set object 66 rect from 4 , 8 to 0.84 , 1 fc rgb "cyan" fillstyle solid
set object 67 rect from 2 , 4 to 0.84 , 1 fc rgb "cyan" fillstyle solid
set object 68 rect from 1 , 2 to 0.84 , 1 fc rgb "cyan" fillstyle solid
set object 69 rect from 0.5 , 1 to 0.84 , 1 fc rgb "cyan" fillstyle solid
set object 70 rect from 0.25 , 0.5 to 0.84 , 1 fc rgb "cyan" fillstyle solid
set object 71 rect from 0.18 , 0.25 to 0.84 , 1 fc rgb "cyan" fillstyle solid
set object 72 rect from 0.15 , 0.18 to 0.84 , 1 fc rgb "cyan" fillstyle solid
set object 73 rect from 20 , 100 to 0.74 , 0.84 fc rgb "cyan" fillstyle solid
set object 74 rect from 8 , 20 to 0.74 , 0.84 fc rgb "cyan" fillstyle solid
set object 75 rect from 4 , 8 to 0.74 , 0.84 fc rgb "cyan" fillstyle solid
set object 76 rect from 2 , 4 to 0.74 , 0.84 fc rgb "cyan" fillstyle solid
set object 77 rect from 1 , 2 to 0.74 , 0.84 fc rgb "cyan" fillstyle solid
set object 78 rect from 0.5 , 1 to 0.74 , 0.84 fc rgb "cyan" fillstyle solid
set object 79 rect from 0.25 , 0.5 to 0.74 , 0.84 fc rgb "cyan" fillstyle solid
set object 80 rect from 0.18 , 0.25 to 0.74 , 0.84 fc rgb "cyan" fillstyle solid
set object 81 rect from 0.15 , 0.18 to 0.74 , 0.84 fc rgb "cyan" fillstyle solid
set object 82 rect from 20 , 100 to 0.65 , 0.74 fc rgb "cyan" fillstyle solid
set object 83 rect from 8 , 20 to 0.65 , 0.74 fc rgb "cyan" fillstyle solid
set object 84 rect from 4 , 8 to 0.65 , 0.74 fc rgb "cyan" fillstyle solid
set object 85 rect from 2 , 4 to 0.65 , 0.74 fc rgb "cyan" fillstyle solid
set object 86 rect from 1 , 2 to 0.65 , 0.74 fc rgb "cyan" fillstyle solid
set object 87 rect from 0.5 , 1 to 0.65 , 0.74 fc rgb "cyan" fillstyle solid
set object 88 rect from 0.25 , 0.5 to 0.65 , 0.74 fc rgb "cyan" fillstyle solid
set object 89 rect from 0.18 , 0.25 to 0.65 , 0.74 fc rgb "cyan" fillstyle solid
set object 90 rect from 0.15 , 0.18 to 0.65 , 0.74 fc rgb "cyan" fillstyle solid
set object 91 rect from 20 , 100 to 0.64 , 0.65 fc rgb "cyan" fillstyle solid
set object 92 rect from 8 , 20 to 0.64 , 0.65 fc rgb "cyan" fillstyle solid
set object 93 rect from 4 , 8 to 0.64 , 0.65 fc rgb "cyan" fillstyle solid
set object 94 rect from 2 , 4 to 0.64 , 0.65 fc rgb "cyan" fillstyle solid
set object 95 rect from 1 , 2 to 0.64 , 0.65 fc rgb "cyan" fillstyle solid
set object 96 rect from 0.5 , 1 to 0.64 , 0.65 fc rgb "cyan" fillstyle solid
set object 97 rect from 0.25 , 0.5 to 0.64 , 0.65 fc rgb "cyan" fillstyle solid
set object 98 rect from 0.18 , 0.25 to 0.64 , 0.65 fc rgb "cyan" fillstyle solid
set object 99 rect from 0.15 , 0.18 to 0.64 , 0.65 fc rgb "cyan" fillstyle solid
set object 100 rect from 20 , 100 to 0.61 , 0.64 fc rgb "cyan" fillstyle solid
set object 101 rect from 8 , 20 to 0.61 , 0.64 fc rgb "cyan" fillstyle solid
set object 102 rect from 4 , 8 to 0.61 , 0.64 fc rgb "cyan" fillstyle solid
set object 103 rect from 2 , 4 to 0.61 , 0.64 fc rgb "cyan" fillstyle solid
set object 104 rect from 1 , 2 to 0.61 , 0.64 fc rgb "cyan" fillstyle solid
set object 105 rect from 0.5 , 1 to 0.61 , 0.64 fc rgb "cyan" fillstyle solid
set object 106 rect from 0.25 , 0.5 to 0.61 , 0.64 fc rgb "cyan" fillstyle solid
set object 107 rect from 0.18 , 0.25 to 0.61 , 0.64 fc rgb "cyan" fillstyle solid
set object 108 rect from 0.15 , 0.18 to 0.61 , 0.64 fc rgb "cyan" fillstyle solid
set object 109 rect from 20 , 100 to 0.6 , 0.61 fc rgb "cyan" fillstyle solid
set object 110 rect from 8 , 20 to 0.6 , 0.61 fc rgb "cyan" fillstyle solid
set object 111 rect from 4 , 8 to 0.6 , 0.61 fc rgb "cyan" fillstyle solid
set object 112 rect from 2 , 4 to 0.6 , 0.61 fc rgb "cyan" fillstyle solid
set object 113 rect from 1 , 2 to 0.6 , 0.61 fc rgb "cyan" fillstyle solid
set object 114 rect from 0.5 , 1 to 0.6 , 0.61 fc rgb "cyan" fillstyle solid
set object 115 rect from 0.25 , 0.5 to 0.6 , 0.61 fc rgb "cyan" fillstyle solid
set object 116 rect from 0.18 , 0.25 to 0.6 , 0.61 fc rgb "cyan" fillstyle solid
set object 117 rect from 0.15 , 0.18 to 0.6 , 0.61 fc rgb "cyan" fillstyle solid
set object 118 rect from 20 , 100 to 0.58 , 0.6 fc rgb "cyan" fillstyle solid
set object 119 rect from 8 , 20 to 0.58 , 0.6 fc rgb "cyan" fillstyle solid
set object 120 rect from 4 , 8 to 0.58 , 0.6 fc rgb "cyan" fillstyle solid
set object 121 rect from 2 , 4 to 0.58 , 0.6 fc rgb "cyan" fillstyle solid
set object 122 rect from 1 , 2 to 0.58 , 0.6 fc rgb "cyan" fillstyle solid
set object 123 rect from 0.5 , 1 to 0.58 , 0.6 fc rgb "cyan" fillstyle solid
set object 124 rect from 0.25 , 0.5 to 0.58 , 0.6 fc rgb "cyan" fillstyle solid
set object 125 rect from 0.18 , 0.25 to 0.58 , 0.6 fc rgb "cyan" fillstyle solid
set object 126 rect from 0.15 , 0.18 to 0.58 , 0.6 fc rgb "cyan" fillstyle solid
set object 127 rect from 20 , 100 to 0.55 , 0.58 fc rgb "cyan" fillstyle solid
set object 128 rect from 8 , 20 to 0.55 , 0.58 fc rgb "cyan" fillstyle solid
set object 129 rect from 4 , 8 to 0.55 , 0.58 fc rgb "cyan" fillstyle solid
set object 130 rect from 2 , 4 to 0.55 , 0.58 fc rgb "cyan" fillstyle solid
set object 131 rect from 1 , 2 to 0.55 , 0.58 fc rgb "cyan" fillstyle solid
set object 132 rect from 0.5 , 1 to 0.55 , 0.58 fc rgb "cyan" fillstyle solid
set object 133 rect from 0.25 , 0.5 to 0.55 , 0.58 fc rgb "cyan" fillstyle solid
set object 134 rect from 0.18 , 0.25 to 0.55 , 0.58 fc rgb "cyan" fillstyle solid
set object 135 rect from 0.15 , 0.18 to 0.55 , 0.58 fc rgb "cyan" fillstyle solid
set object 136 rect from 20 , 100 to 0.54 , 0.55 fc rgb "cyan" fillstyle solid
set object 137 rect from 8 , 20 to 0.54 , 0.55 fc rgb "cyan" fillstyle solid
set object 138 rect from 4 , 8 to 0.54 , 0.55 fc rgb "cyan" fillstyle solid
set object 139 rect from 2 , 4 to 0.54 , 0.55 fc rgb "cyan" fillstyle solid
set object 140 rect from 1 , 2 to 0.54 , 0.55 fc rgb "cyan" fillstyle solid
set object 141 rect from 0.5 , 1 to 0.54 , 0.55 fc rgb "cyan" fillstyle solid
set object 142 rect from 0.25 , 0.5 to 0.54 , 0.55 fc rgb "cyan" fillstyle solid
set object 143 rect from 0.18 , 0.25 to 0.54 , 0.55 fc rgb "cyan" fillstyle solid
set object 144 rect from 0.15 , 0.18 to 0.54 , 0.55 fc rgb "cyan" fillstyle solid
set object 145 rect from 20 , 100 to 0.52 , 0.54 fc rgb "cyan" fillstyle solid
set object 146 rect from 8 , 20 to 0.52 , 0.54 fc rgb "cyan" fillstyle solid
set object 147 rect from 4 , 8 to 0.52 , 0.54 fc rgb "cyan" fillstyle solid
set object 148 rect from 2 , 4 to 0.52 , 0.54 fc rgb "cyan" fillstyle solid
set object 149 rect from 1 , 2 to 0.52 , 0.54 fc rgb "cyan" fillstyle solid
set object 150 rect from 0.5 , 1 to 0.52 , 0.54 fc rgb "cyan" fillstyle solid
set object 151 rect from 0.25 , 0.5 to 0.52 , 0.54 fc rgb "cyan" fillstyle solid
set object 152 rect from 0.18 , 0.25 to 0.52 , 0.54 fc rgb "cyan" fillstyle solid
set object 153 rect from 0.15 , 0.18 to 0.52 , 0.54 fc rgb "cyan" fillstyle solid
set object 154 rect from 20 , 100 to 0.42 , 0.52 fc rgb "cyan" fillstyle solid
set object 155 rect from 8 , 20 to 0.42 , 0.52 fc rgb "cyan" fillstyle solid
set object 156 rect from 4 , 8 to 0.42 , 0.52 fc rgb "cyan" fillstyle solid
set object 157 rect from 2 , 4 to 0.42 , 0.52 fc rgb "cyan" fillstyle solid
set object 158 rect from 1 , 2 to 0.42 , 0.52 fc rgb "cyan" fillstyle solid
set object 159 rect from 0.5 , 1 to 0.42 , 0.52 fc rgb "cyan" fillstyle solid
set object 160 rect from 0.25 , 0.5 to 0.42 , 0.52 fc rgb "cyan" fillstyle solid
set object 161 rect from 0.18 , 0.25 to 0.42 , 0.52 fc rgb "cyan" fillstyle solid
set object 162 rect from 0.15 , 0.18 to 0.42 , 0.52 fc rgb "cyan" fillstyle solid
set object 163 rect from 20 , 100 to 0.39 , 0.42 fc rgb "cyan" fillstyle solid
set object 164 rect from 8 , 20 to 0.39 , 0.42 fc rgb "cyan" fillstyle solid
set object 165 rect from 4 , 8 to 0.39 , 0.42 fc rgb "cyan" fillstyle solid
set object 166 rect from 2 , 4 to 0.39 , 0.42 fc rgb "cyan" fillstyle solid
set object 167 rect from 1 , 2 to 0.39 , 0.42 fc rgb "cyan" fillstyle solid
set object 168 rect from 0.5 , 1 to 0.39 , 0.42 fc rgb "cyan" fillstyle solid
set object 169 rect from 0.25 , 0.5 to 0.39 , 0.42 fc rgb "cyan" fillstyle solid
set object 170 rect from 0.18 , 0.25 to 0.39 , 0.42 fc rgb "cyan" fillstyle solid
set object 171 rect from 0.15 , 0.18 to 0.39 , 0.42 fc rgb "cyan" fillstyle solid
set object 172 rect from 20 , 100 to 0.36 , 0.39 fc rgb "cyan" fillstyle solid
set object 173 rect from 8 , 20 to 0.36 , 0.39 fc rgb "cyan" fillstyle solid
set object 174 rect from 4 , 8 to 0.36 , 0.39 fc rgb "cyan" fillstyle solid
set object 175 rect from 2 , 4 to 0.36 , 0.39 fc rgb "cyan" fillstyle solid
set object 176 rect from 1 , 2 to 0.36 , 0.39 fc rgb "cyan" fillstyle solid
set object 177 rect from 0.5 , 1 to 0.36 , 0.39 fc rgb "cyan" fillstyle solid
set object 178 rect from 0.25 , 0.5 to 0.36 , 0.39 fc rgb "cyan" fillstyle solid
set object 179 rect from 0.18 , 0.25 to 0.36 , 0.39 fc rgb "cyan" fillstyle solid
set object 180 rect from 0.15 , 0.18 to 0.36 , 0.39 fc rgb "cyan" fillstyle solid
